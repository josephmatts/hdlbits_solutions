module simple_wire
(
    input  in, 
    output out
);

    assign out = in;

endmodule