module gnd 
(
    output out
);
	assign out = 0;
endmodule
